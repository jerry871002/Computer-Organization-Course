// 0610780

//Subject:     CO project 2 - Sign extend
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:
//----------------------------------------------
//Date:
//----------------------------------------------
//Description:
//--------------------------------------------------------------------------------

module Sign_Extend(
    data_i,
    data_o
    );

//I/O ports
input   [16-1:0] data_i;
output  [32-1:0] data_o;

//Internal Signals
reg     [32-1:0] data_o;

//Sign extended
always @ ( * ) begin
    if (data_i[15]) begin
        data_o <= { 16'hffff, data_i[15:0] };
    end else begin
        data_o <= { 16'h0000, data_i[15:0] };
    end
end

endmodule
