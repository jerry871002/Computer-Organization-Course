//Subject:     CO project 2 - Decoder
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      Luke
//----------------------------------------------
//Date:        2010/8/16
//----------------------------------------------
//Description:
//--------------------------------------------------------------------------------

module Decoder(
    instr_op_i,
	RegWrite_o,
	ALU_op_o,
	ALUSrc_o,
	RegDst_o,
	Branch_o,
    Jump_o,
    MemRead_o,
    MemWrite_o,
    MemtoReg_o
	);

//I/O ports
input  [6-1:0] instr_op_i;

output         RegWrite_o;
output [3-1:0] ALU_op_o;
output         ALUSrc_o;
output         RegDst_o;
output         Branch_o;
output         Jump_o;
output         MemRead_o;
output         MemWrite_o;
output         MemtoReg_o;

//Internal Signals
reg    [3-1:0] ALU_op_o;
reg            ALUSrc_o;
reg            RegWrite_o;
reg            RegDst_o;
reg            Branch_o;
reg            Jump_o;
reg            MemRead_o;
reg            MemWrite_o;
reg            MemtoReg_o;

//Parameter

//Main function
always @ ( * ) begin
    case(instr_op_i)
        // jal
        6'b000011: begin
            RegWrite_o <= 1'b1;
            ALU_op_o <= 3'b011;
            RegDst_o <= 1'bx;
            Branch_o <= 1'b0;
            Jump_o <= 1'b1;
            MemRead_o <= 1'b0;
            MemWrite_o <= 1'b0;
            MemtoReg_o <= 1'bx;
        end
        // lw
        6'b100011: begin
            RegWrite_o <= 1'b1;
            ALU_op_o <= 3'b110;
            RegDst_o <= 1'b0;
            Branch_o <= 1'b0;
            Jump_o <= 1'b0;
            MemRead_o <= 1'b1;
            MemWrite_o <= 1'b0;
            MemtoReg_o <= 1'b1;
        end
        // sw
        6'b101011: begin
            RegWrite_o <= 1'b0;
            ALU_op_o <= 3'b110;
            RegDst_o <= 1'b0;
            Branch_o <= 1'b0;
            Jump_o <= 1'b0;
            MemRead_o <= 1'b0;
            MemWrite_o <= 1'b1;
            MemtoReg_o <= 1'b0;
        end
        // jump
        6'b000010: begin
            RegWrite_o <= 1'b0;
            ALU_op_o <= 3'b011;
            RegDst_o <= 1'b1;
            Branch_o <= 1'b0;
            Jump_o <= 1'b1;
            MemRead_o <= 1'b0;
            MemWrite_o <= 1'b0;
            MemtoReg_o <= 1'b0;
        end
        // beq
        6'b000100: begin
            RegWrite_o <= 1'b0;
            ALU_op_o <= 3'b011;
            RegDst_o <= 1'b1;
            Branch_o <= 1'b1;
            Jump_o <= 1'b0;
            MemRead_o <= 1'b0;
            MemWrite_o <= 1'b0;
            MemtoReg_o <= 1'b0;
        end
        // addi
        6'b001000: begin
            RegWrite_o <= 1'b1;
            ALU_op_o <= 3'b110;
            RegDst_o <= 1'b0;
            Branch_o <= 1'b0;
            Jump_o <= 1'b0;
            MemRead_o <= 1'b0;
            MemWrite_o <= 1'b0;
            MemtoReg_o <= 1'b0;
        end
        // R-type
        default: begin
            RegWrite_o <= 1'b1;
            ALU_op_o <= 3'b000;
            RegDst_o <= 1'b1;
            Branch_o <= 1'b0;
            Jump_o <= 1'b0;
            MemRead_o <= 1'b0;
            MemWrite_o <= 1'b0;
            MemtoReg_o <= 1'b0;
        end
    endcase

    ALUSrc_o <= instr_op_i[3] | instr_op_i[5];

end

endmodule
